`include "cpu/pipelineInterfaces.sv"
module ID (
    input      clk,
    input      rst,
    IController.ID i_controller,
    IIF_ID.ID i_if_id,
    input [37:0]WB_BACK,
    input [37:0]MEM_BACK,
    input [31:2]CP0_EPC,
    output reg[15:0]o_EX_CTRL,
    output reg o_MEM_CTRL,
    output reg [4:0] o_WB_CTRL,
    output reg[157:0] o_EX_DATA,
);  
    wire [2:0]branchType;
    assign {NPCFromEPC,ExlSet,jmp,NPCFromGPR,branchType,extop,exsign}=i_controller.ID_CTRL;
    assign o_uncertainJump=NPCFromGPR||(branchType!=0);
    wire [31:2] PCP1;
    wire [31:0] instr;
    assign {PCP1,instr}=i_if_id.ID_DATA;
    assign i_controller.ID_instr=instr;
    wire [31:0] WB_Wd;
    wire [4:0] WB_rw;
    assign {WB_regWrite,WB_Wd,WB_rw}=WB_BACK;

    wire [31:0]rd1,rd2,EXTB;

    GPR GPR(
        .clk(clk),  //for WB befor ID
        .reset(rst),
        .rs(instr[25:21]),
        .rt(instr[20:16]),
        .rw(WB_rw),
        .regWrite(WB_regWrite),
        .Wd(WB_Wd),
        .rd1(rd1),
        .rd2(rd2) 
    );
 
    EXT EXT(
        .A(instr[15:0]),
        .extop(extop),
        .exsign(exsign),
        .B(EXTB)
    );
    // outports wire
    wire [31:0] 	f_rd1;
    wire [31:0] 	f_rd2;
    
    FORWARD u_ID_FORWARD(
        .MEM_BACK 	( MEM_BACK  ),
        .WB_BACK  	( WB_BACK   ),
        .USE_MEM_BACK(1'b1),
        .USE_WB_BACK(1'b1),
        .rs       	( instr[25:21]       ),
        .rt       	( instr[20:16]        ),
        .rd1      	( rd1       ),
        .rd2      	( rd2       ),
        .f_rd1    	( f_rd1     ),
        .f_rd2    	( f_rd2     )
    );
    // outports wire
    wire       	branchAvail;
    
    BRANCH u_BRANCH(
        .rd1          	( f_rd1           ),
        .rd2        	( f_rd2         ),
        .branchType  	( branchType   ),
        .branchAvail 	( branchAvail  )
    );
    
    jpc jpc (
        .PC(PCP1),
        .branchAvail(branchAvail), 
        .jmp(jmp),
        .offset(instr[15:0]),
        .instr_index(instr[25:0]),
        .reg_index(f_rd1),
        .NPCFromGPR(NPCFromGPR),
        .goExceptionHandler(ExlSet),
        .NPCFromEPC(NPCFromEPC),
        .EPC(CP0_EPC),
        .JPC(i_if_id.JPC)
    );

    assign i_if_id.jpcAvail=ExlSet|NPCFromEPC||NPCFromGPR||jmp||branchAvail;
    initial begin
        o_EX_DATA<=0;
        o_EX_CTRL<=0;
        o_MEM_CTRL<=0;
        o_WB_CTRL<=0;
    end
    always @(posedge clk) begin
        if(i_controller.ID_FLUSH) begin
            //o_EX_DATA<=0;
            o_EX_CTRL<=0;
            o_MEM_CTRL<=0;
            o_WB_CTRL<=0;
        end
        else begin
            o_EX_DATA<={PCP1,instr,f_rd1,f_rd2,EXTB};
            o_EX_CTRL<=i_controller.EX_CTRL;
            o_MEM_CTRL<=i_controller.MEM_CTRL;
            o_WB_CTRL<=i_controller.WB_CTRL;
        end
    end
endmodule //ID